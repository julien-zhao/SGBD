�� sr java.util.ArrayListx����a� I sizexp   w   sr RelationInfo        L headerPageIdt LPageId;L nomRelationt Ljava/lang/String;L tabInfot Ljava/util/List;xpsr PageId        I fileIdxI pageIdxxp        t Ssq ~     w   sr ColInfo        L colonneq ~ L typeq ~ xpt C1t INTEGERsq ~ t C2t REALsq ~ t C3t INTEGERsq ~ t C4t INTEGERsq ~ t C5t INTEGERxx