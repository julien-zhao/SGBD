�� sr java.util.ArrayListx����a� I sizexp   w   sr RelationInfo        L headerPageIdt LPageId;L nomRelationt Ljava/lang/String;L tabInfot Ljava/util/List;xppt RelationNonVidesq ~     w   sr ColInfo        L colonneq ~ L typeq ~ xpt Nomt VARCHAR(10)sq ~ 	t Prenomt VARCHAR(12)sq ~ 	t Aget INTEGERsq ~ 	t NoteEXt REALxsq ~ pt RelationQuiEstVidesq ~      w    xx