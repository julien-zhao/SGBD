�� sr java.util.ArrayListx����a� I sizexp   w   sr RelationInfo        L headerPageIdt LPageId;L nomRelationt Ljava/lang/String;L tabInfot Ljava/util/List;xpsr PageId        I fileIdxI pageIdxxp        t RelationNonVidesq ~     w   sr ColInfo        L colonneq ~ L typeq ~ xpt Nomt VARCHAR(10)sq ~ t Prenomt VARCHAR(12)sq ~ t Aget INTEGERsq ~ t NoteEXt REALxsq ~ sq ~         t RelationQuiEstVidesq ~      w    xx