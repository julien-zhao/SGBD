�� sr java.util.ArrayListx����a� I sizexp   w   {sr  java.io.NotSerializableException(Vx �5  xr java.io.ObjectStreamExceptiond��k�9��  xr java.io.IOExceptionl�sde%�  xr java.lang.Exception��>;�  xr java.lang.Throwable��5'9w�� L causet Ljava/lang/Throwable;L detailMessaget Ljava/lang/String;[ 
stackTracet [Ljava/lang/StackTraceElement;L suppressedExceptionst Ljava/util/List;xpq ~ 	t RelationInfour [Ljava.lang.StackTraceElement;F*<<�"9  xp   sr java.lang.StackTraceElementa	Ś&6݅ B formatI 
lineNumberL classLoaderNameq ~ L declaringClassq ~ L fileNameq ~ L 
methodNameq ~ L 
moduleNameq ~ L moduleVersionq ~ xp  �pt java.io.ObjectOutputStreamt ObjectOutputStream.javat writeObject0t 	java.baset 17.0.3sq ~   bpq ~ q ~ t writeObjectq ~ q ~ sq ~   bpt java.util.ArrayListt ArrayList.javaq ~ q ~ q ~ sq ~ ����pt -jdk.internal.reflect.NativeMethodAccessorImplt NativeMethodAccessorImpl.javat invoke0q ~ q ~ sq ~    Mpq ~ q ~ t invokeq ~ q ~ sq ~    +pt 1jdk.internal.reflect.DelegatingMethodAccessorImplt !DelegatingMethodAccessorImpl.javaq ~ q ~ q ~ sq ~   8pt java.lang.reflect.Methodt Method.javaq ~ q ~ q ~ sq ~   �pt java.io.ObjectStreamClasst ObjectStreamClass.javat invokeWriteObjectq ~ q ~ sq ~   �pq ~ q ~ t writeSerialDataq ~ q ~ sq ~   �pq ~ q ~ t writeOrdinaryObjectq ~ q ~ sq ~   �pq ~ q ~ q ~ q ~ q ~ sq ~   bpq ~ q ~ q ~ q ~ q ~ sq ~    #t appt Catalogt Catalog.javat Finishppsq ~    q ~ 0t CatalogTestt CatalogTest.javat mainppsr java.util.Collections$EmptyListz��<���  xpx